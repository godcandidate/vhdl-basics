----------------------------------------------------------------------------------
-- Company: 
-- Engineer:  Eddie
-- 
-- Create Date:    20:59:25 07/27/2023 
-- Design Name: 	Eddie
-- Module Name:    and_gate - Dataflow 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity and_gate is
end and_gate;

architecture Dataflow of and_gate is

begin


end Dataflow;

